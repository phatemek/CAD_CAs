module Not(x, nx);input x;output nx;C2 myc2(1'b1, 1'b1, 1'b1, 1'b0, x, x, x, x, nx);endmodule
