module reg10bit(A, clk, rst, out);input clk, rst;input [9:0] A;output [9:0] out;wire b9, b8, b7, b6, b5, b4, b3, b2, b1, b0;S2 reg9(A[9], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rst, clk, b9);S2 reg8(A[8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b8);S2 reg7(A[7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b7);S2 reg6(A[6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b6);S2 reg5(A[5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rst, clk, b5);S2 reg4(A[4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b4);S2 reg3(A[3], 01'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b3);S2 reg2(A[2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b2);S2 reg1(A[1], 01'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b1);S2 reg0(A[0], 01'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  rst, clk, b0);assign out = {b9, b8, b7, b6, b5, b4, b3, b2, b1, b0};endmodule
