module Co(a, b, c, out);input a, b, c;output out;C2 myc2(1'b0, c, c, 1'b1, a, b, a, b, out);endmodule
