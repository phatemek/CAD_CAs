module Actfun(A, out);input [11:0] A;output [4:0] out;wire lb;wire[11:0] B;assign lb = A[11];C2 c0(A[11], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[11]);C2 c1(A[10], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[10]);C2 c2(A[9], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[9]);C2 c3(A[8], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[8]);C2 c4(A[7], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[7]);C2 c5(A[6], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[6]);C2 c6(A[5], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[5]);C2 c7(A[4], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[4]);C2 c8(A[3], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[3]);C2 c9(A[2], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[2]);C2 c10(A[1], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[1]);C2 c11(A[0], 1'b0, 1'b0, 1'b0, lb, lb, lb, lb, B[0]);assign out = {B[11], B[6:3]};endmodule
