module Adder(a, b, out);
	input [8:0] a, b;
	output [8:0] out;
	assign out = a + b;
endmodule	
