module And5bit(a, b, res);input [4:0] a, b;output [4:0] res;C2 myc21(1'b0, 1'b0, 1'b0, 1'b1, a[4], b[4], a[4], b[4], res[4]);C2 myc22(1'b0, 1'b0, 1'b0, 1'b1, a[3], b[3], a[3], b[3], res[3]);C2 myc23(1'b0, 1'b0, 1'b0, 1'b1, a[2], b[2], a[2], b[2], res[2]);C2 myc24(1'b0, 1'b0, 1'b0, 1'b1, a[1], b[1], a[1], b[1], res[1]);C2 myc25(1'b0, 1'b0, 1'b0, 1'b1, a[0], b[0], a[0], b[0], res[0]);endmodule
