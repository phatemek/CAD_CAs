module Or1bit(a0, a1, a2, a3, a4, a5, out);input a0, a1, a2, a3, a4, a5;output out;wire w1, w2, w3, w4;C2 myc21(1'b0, 1'b1, 1'b1, 1'b1, a0, a1, a0, a1, w1);C2 myc22(1'b0, 1'b1, 1'b1, 1'b1, a2, a3, a2, a3, w2);C2 myc23(1'b0, 1'b1, 1'b1, 1'b1, a4, a5, a4, a5, w3);C2 myc24(1'b0, 1'b1, 1'b1, 1'b1, w1, w2, w1, w2, w4);C2 myc25(1'b0, 1'b1, 1'b1, 1'b1, w4, w3, w4, w3, out);endmodule
